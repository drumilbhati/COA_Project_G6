module ALU(clk, Reset, Imm7, Op1, Op2, OpCode, ALU_Save, ZFlag_Save, CFlag_Save);

endmodule